spice test 4-diode bridge circuit + 1 diode
* 4-diode circuit under 2-tone excitation
* "t" transmission line included  
* large LO signal
*
*
*
*


vs  1 0  ac 1v sin (0 21.21 100Meg 0 0) 
+              distof1 15 

*t1  1 0 2 0 z0=50 f=100MEG nl=0.5 
rr 1 2 2

d1 2 3 sd
d2 4 2 sd
d3 5 3 sd
d4 4 5 sd

rg 5 0 2

d5 6 7  sd 
d6 6 7  sd
rs1 2 6 2 
rs2 7 0 2

rl  3 4  1k


.model sd d is=1e-9 tt=0 m=0.5

* .ac dec 5 10 10k 
.tran 0.2n 500n 0 0.2n

.hb f1=100e6 f2=0 
+ 0 0 1 0 2 0 3 0 4 0 5 0  
+ 6 0 7 0 8 0 9 0 10 0 
+ 11 0 12 0 13 0 14 0 15 0 
+ 16 0 17 0 18 0 19 0  

.hb_options epsiw=1.e-6 epssol=1.e-12 epsdu=1.e-9 limit=50


.end
